module flash_read(

    input               clk         ,
    input               rst_n       ,
    
    //key
    input               rd_id       ,
    input               rd_data     ,
    
    input   [23:0]      rd_addr     ,//flash读地址

    //spi_master
    output              trans_req   ,
    output  [7:0]       tx_dout     ,
    input   [7:0]       rx_din      ,
    input               trans_done  ,

    //output
    output  [47:0]      dout        ,
    output  [5:0]       dout_mask   ,
    output              dout_vld    
);

/*********  工程注释        ****************

M25P16 Flash读控制器，实现读数据和读存储器的ID。

**********  注释结束    ****************/

//状态机参数定义
    localparam  IDLE = 4'b0001,
                RDID = 4'b0010,//读器件ID
                RDDA = 4'b0100,//读数据字节
                DONE = 4'b1000;
//Flash命令参数定义
    localparam  CMD_RDID = 8'h9F,
                CMD_RDDA = 8'h03;

//信号定义

    reg     [3:0]       state_c     ;
    reg     [3:0]       state_n     ;

    reg     [3:0]       cnt_byte    ;
    wire                add_cnt_byte;
    wire                end_cnt_byte;
    reg     [3:0]       byte_num    ;

    reg     [7:0]       tx_data     ;
    reg                 tx_req      ;
    
    reg                 flag        ;//读数据、读ID标志

    wire                idle2rdid   ; 
    wire                rdid2done   ; 
    wire                idle2rdda   ; 
    wire                rdda2done   ; 
    wire                done2idle   ; 
    
    reg     [31:0]      rx_data	/* synthesis keep */;//串并转换寄存器
    reg     [47:0]      data        ;
    reg     [5:0]       data_mask   ;
    reg                 data_vld    ;

//状态机
    
    always @(posedge clk or negedge rst_n) begin 
        if (rst_n==0) begin
            state_c <= IDLE ;
        end
        else begin
            state_c <= state_n;
       end
    end
    
    always @(*) begin 
        case(state_c)  
            IDLE :begin
                if(idle2rdid)
                    state_n = RDID ;
                else if(idle2rdda)
                    state_n = RDDA ;
                else 
                    state_n = state_c ;
            end
            RDID :begin
                if(rdid2done)
                    state_n = DONE ;
                else 
                    state_n = state_c ;
            end
            RDDA :begin
                if(rdda2done)
                    state_n = DONE ;
                else 
                    state_n = state_c ;
            end
            DONE :begin
                if(done2idle)
                    state_n = IDLE ;
                else 
                    state_n = state_c ;
            end
            default : state_n = IDLE ;
        endcase
    end
    
    assign idle2rdid = state_c==IDLE && (rd_id  );
    assign rdid2done = state_c==RDID && (end_cnt_byte);
    assign idle2rdda = state_c==IDLE && (rd_data);
    assign rdda2done = state_c==RDDA && (end_cnt_byte);
    assign done2idle = state_c==DONE && (1'b1);
    
    always @(posedge clk or negedge rst_n) begin 
        if (rst_n==0) begin
            cnt_byte <= 0; 
        end
        else if(add_cnt_byte) begin
            if(end_cnt_byte)
                cnt_byte <= 0; 
            else
                cnt_byte <= cnt_byte+1 ;
       end
    end
    assign add_cnt_byte = (state_c != IDLE && trans_done);
    assign end_cnt_byte = add_cnt_byte  && cnt_byte == (byte_num)-1 ;
        
    always  @(*)begin
        if(state_c == RDID)
            byte_num = 4;
        else  
            byte_num = 8;   //至少5B CMD + 3 ADDR + X DATA
    end

//输出
    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            tx_req <= 1'b0;
        end
        else if(idle2rdid | idle2rdda)begin
            tx_req <= 1'b1;
        end
        else if(rdid2done | rdda2done)begin
            tx_req <= 1'b0;
        end
    end

    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            tx_data <= 0;
        end
        else if(state_c == RDID)begin
            case(cnt_byte)
                0:tx_data <= CMD_RDID;  
                default:tx_data <= 0; 
            endcase 
        end
        else if(state_c == RDDA)begin
            case(cnt_byte)
                0:tx_data <= CMD_RDDA; 
                1:tx_data <= rd_addr[23:16];
                2:tx_data <= rd_addr[15:8];
                3:tx_data <= rd_addr[7:0];
                default:tx_data <= 0; 
            endcase 
        end
    end

    //rx_data
    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            rx_data <= 0;
        end
        else if(state_c == RDID && trans_done)begin
            rx_data <= {rx_data[23:0],rx_din};
        end
        else if(state_c == RDDA && trans_done)begin
            rx_data <= {rx_data[23:0],rx_din};
        end
    end

    //data  
    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            data <= 0;
        end
        else if(state_c == DONE && ~flag)begin   //读ID
            data <= {4'd0,rx_data[23:20],4'd0,rx_data[19:16],   //2 0
                     4'd0,rx_data[15:12],4'd0,rx_data[11:8],    //2 0
                     4'd0,rx_data[7:4],4'd0,rx_data[3:0]};      //1 5 
        end 
        else if(state_c == DONE && flag)begin //读数据
            data <= {"R","D",16'd0,4'd0,rx_data[7:4],4'd0,rx_data[3:0]};
        end 
    end

    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            data_mask <= 0;
        end
        else if(state_c == DONE && ~flag)begin
            data_mask <= 6'b00_0000;
        end
        else if(state_c == DONE && flag)begin
            data_mask <= 6'b00_1100;
        end
    end

    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            data_vld <= 0;
        end
        else begin
            data_vld <= state_c == DONE; 
        end
    end

    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            flag <= 1'b0;
        end
        else if(idle2rdda)begin
            flag <= 1'b1;
        end
        else if(idle2rdid)begin
            flag <= 1'b0;
        end
    end

//输出
    assign tx_dout =tx_data;
    assign trans_req = tx_req;

    assign dout = data;
    assign dout_mask = data_mask;
    assign dout_vld = data_vld;

endmodule 


